netcdf test_mmr {   // generate date for fixmmr
  dimensions:
	  lon = 4 ;
	  lat = 5 ;
          height = 3;
  variables:
	  float O1(lon, lat,height) ;
	  float O2(lon, lat,height) ;
	  float HE(lon, lat,height) ;
  // global attributes
	  :title = "MMR test data tiegcm";
  data:
   O1 =
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 1.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3;

   O2 =
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 2.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3;

   HE =
    0.3, 3.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3,
    0.3, 0.3, 0.3, 0.3;
  }

